module FIFO(
    input wire i_clk,
    input wire i_rst,
    input wire i_we;
    input wire i_re;
    input wire i_data;
    output wire o_full;
    output wire o_empty;
    output wire o_data;
);
endmodule